--------------------------------------------------------------------
--! \file      ch04_exm04_4.vhd
--! \date      see top of 'Version History'
--! \brief     Example 4.4 of Pedroni 2nd Ed, page 109.
--! \author    Remko Welling (WLGRW) remko.welling@han.nl
--! \copyright HAN TF ELT/ESE Arnhem 
--!
--! Version History:
--! ----------------
--!
--! Nr:    |Date:      |Author: |Remarks:
--! -------|-----------|--------|-----------------------------------
--! 001    |9-12-2019  |WLGRW   |Added architecture switch
--!

--! Function description:
--! ---------------------
--! This implementation is using ATTRIBUTE KEEP to prevent 
--! optimisation of synthesis. As a result the logic is kept and 
--! will introduce delay trough the logic.
--!
--! Assignment:
--! -----------
--! 1- Example 4.4 of Pedroni 2nd Ed, page 109.
--! 2- Compile the code with uncommented KEEP attribute and inspect
--!    Hardware compiled
--! 3- Compile the code with commented KEEP attribute and inspect
--!    Hardware compiled
--! 4- Answer the question: what is changed?


------------------------------------------------------------------
--! Include libraries

------------------------------------------------------------------
--! Add ENTITY



----------------------------------------------------------------
--! Add ARCHITECTURE and IMPLEMENT code 







------------------------------------------------------------------
